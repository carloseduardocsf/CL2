module projeto11_revisao (a, b, c, y, z);

input a, b, c;
output y, z;


endmodule