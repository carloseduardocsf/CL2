module ex10(nen, addr, row_sel);

input nem, addr[2:0];
output row_sel[7:0];




endmodule
