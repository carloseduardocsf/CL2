module projeto08 ();




endmodule